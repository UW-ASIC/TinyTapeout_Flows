magic
tech sky130A
timestamp 1625000000
<< nwell >>
rect 100 100 300 300
<< pwell >>
rect 100 -200 300 0
<< metal1 >>
rect 0 0 50 50
rect 350 0 400 50
rect 175 350 225 400
rect 175 -250 225 -300
<< labels >>
flabel metal1 25 25 25 25 0 FreeSans 200 0 0 0 IN
flabel metal1 375 25 375 25 0 FreeSans 200 0 0 0 OUT
flabel metal1 200 375 200 375 0 FreeSans 200 0 0 0 VDD
flabel metal1 200 -275 200 -275 0 FreeSans 200 0 0 0 VSS
<< end >>
