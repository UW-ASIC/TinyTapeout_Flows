** sch_path: /home/omare/Documents/UWASIC/Template/analog/xschem/schematics/template_tb.sch
**.subckt template_tb
I0 VDD Ib 10u
C1 Vout GND 1p m=1
x1 Vp Vn Vout VDD VSS Ib template
V0 VSS GND 0
V2 VDD GND {vdd}
E1 Vp net2 net1 GND 0.5
E2 Vn net2 net1 GND -0.5
Vdm net1 GND ac 1
Vcm net2 GND {vcm}
**** begin user architecture code


.param vdd=1.8
.param vcm=0.9

.control

    save all

    * operating point
    op

    write template.raw
    set appendwrite

    * run ac simulation
    ac dec 20 1k 100e6

    * measure parameters
    let vout_mag = abs(v(Vout))
    let vout_phase_margin = phase(v(Vout)) * 180/pi + 180
    meas ac A0 find vout_mag at=1k
    meas ac UGF when vout_mag=1 fall=1
    meas ac PM find vout_phase_margin when vout_mag=1

    write template_tb.raw
.endc


?
**** end user architecture code
**.ends
.GLOBAL GND
.end
